

module bcdTo7Seg(
    input [4:0] A,
    output [6:0] sseg
);

assign sseg = 
    (A == 5'b00000) ? 7'b0000001 : // 0
    (A == 5'b00001) ? 7'b1001111 : // 1
    (A == 5'b00010) ? 7'b0010010 : // 2
    (A == 5'b00011) ? 7'b0000110 : // 3
    (A == 5'b00100) ? 7'b1001100 : // 4
    (A == 5'b00101) ? 7'b0100100 : // 5
    (A == 5'b00110) ? 7'b0100000 : // 6
    (A == 5'b00111) ? 7'b0001111 : // 7
    (A == 5'b01000) ? 7'b0000000 : // 8
    (A == 5'b01001) ? 7'b0000100 : // 9
    7'b1111111; // All segments off when input is invalid

endmodule
